-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Nov 12 16:20:55 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maqestados IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z1 : OUT STD_LOGIC;
        Z2 : OUT STD_LOGIC;
        Z3 : OUT STD_LOGIC;
        Z4 : OUT STD_LOGIC
    );
END maqestados;

ARCHITECTURE BEHAVIOR OF maqestados IS
    TYPE type_fstate IS (A1,A2,A3,A4,B2,B3,B4,B5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN
            fstate <= A1;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,x)
    BEGIN
        Z1 <= '0';
        Z2 <= '0';
        Z3 <= '0';
        Z4 <= '0';
        CASE fstate IS
            WHEN A1 =>
                IF ((x = '0')) THEN
                    reg_fstate <= A2;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= B2;
                END IF;

                Z1 <= '0';

                Z4 <= '0';

                Z2 <= '0';

                Z3 <= '0';
            WHEN A2 =>
                reg_fstate <= A3;

                Z1 <= '0';

                Z4 <= '0';

                Z2 <= '1';

                Z3 <= '1';
            WHEN A3 =>
                IF ((x = '0')) THEN
                    reg_fstate <= A4;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= B4;
                END IF;

                Z1 <= '1';

                Z4 <= '1';

                Z2 <= '1';

                Z3 <= '1';
            WHEN A4 =>
                reg_fstate <= A1;

                Z1 <= '1';

                Z4 <= '1';

                Z2 <= '0';

                Z3 <= '0';
            WHEN B2 =>
                reg_fstate <= B3;

                Z1 <= '1';

                Z4 <= '0';

                Z2 <= '0';

                Z3 <= '0';
            WHEN B3 =>
                reg_fstate <= B4;

                Z1 <= '1';

                Z4 <= '0';

                Z2 <= '1';

                Z3 <= '0';
            WHEN B4 =>
                IF ((x = '0')) THEN
                    reg_fstate <= A3;
                ELSIF ((x = '1')) THEN
                    reg_fstate <= B5;
                END IF;

                Z1 <= '1';

                Z4 <= '1';

                Z2 <= '1';

                Z3 <= '1';
            WHEN B5 =>
                reg_fstate <= A1;

                Z1 <= '1';

                Z4 <= '0';

                Z2 <= '1';

                Z3 <= '1';
            WHEN OTHERS => 
                Z1 <= 'X';
                Z2 <= 'X';
                Z3 <= 'X';
                Z4 <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
