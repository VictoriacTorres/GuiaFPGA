library verilog;
use verilog.vl_types.all;
entity ej_combinaiconal_vlg_vec_tst is
end ej_combinaiconal_vlg_vec_tst;
